
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;
use IEEE.FIXED_PKG.all;

PACKAGE cordic_pkg IS

    TYPE t_tan_ceoffs_real IS ARRAY(integer RANGE <>) OF real;
    TYPE t_tan_ceoffs_sfixed IS ARRAY(integer RANGE <>) OF sfixed(7 downto -24);
    
    CONSTANT C_K : sfixed(7 downto -24) := to_sfixed(0.6072529350088814, 7, -24);
    
    CONSTANT C_TANGENT_TABLE_REAL: t_tan_ceoffs_real(0 to 31) := (
        0.7853981633974483,
        0.4636476090008061,
        0.24497866312686414,
        0.12435499454676144,
        0.06241880999595735,
        0.031239833430268277,
        0.015623728620476831,
        0.007812341060101111,
        0.0039062301319669718,
        0.0019531225164788188,
        0.0009765621895593195,
        0.0004882812111948983,
        0.00024414062014936177,
        0.00012207031189367021,
        6.103515617420877e-05,
        3.0517578115526096e-05,
        1.5258789061315762e-05,
        7.62939453110197e-06,
        3.814697265606496e-06,
        1.907348632810187e-06,
        9.536743164059608e-07,
        4.7683715820308884e-07,
        2.3841857910155797e-07,
        1.1920928955078068e-07,
        5.960464477539055e-08,
        2.9802322387695303e-08,
        1.4901161193847655e-08,
        7.450580596923828e-09,
        3.725290298461914e-09,
        1.862645149230957e-09,
        9.313225746154785e-10,
        4.656612873077393e-10
    );

    CONSTANT C_TANGENT_TABLE_SFIXED: t_tan_ceoffs_sfixed(0 to 31) := (
        to_sfixed(0.7853981633974483, 7, -24),
        to_sfixed(0.4636476090008061, 7, -24),
        to_sfixed(0.24497866312686414, 7, -24),
        to_sfixed(0.12435499454676144, 7, -24),
        to_sfixed(0.06241880999595735, 7, -24),
        to_sfixed(0.031239833430268277, 7, -24),
        to_sfixed(0.015623728620476831, 7, -24),
        to_sfixed(0.007812341060101111, 7, -24),
        to_sfixed(0.0039062301319669718, 7, -24),
        to_sfixed(0.0019531225164788188, 7, -24),
        to_sfixed(0.0009765621895593195, 7, -24),
        to_sfixed(0.0004882812111948983, 7, -24),
        to_sfixed(0.00024414062014936177, 7, -24),
        to_sfixed(0.00012207031189367021, 7, -24),
        to_sfixed(6.103515617420877e-05, 7, -24),
        to_sfixed(3.0517578115526096e-05, 7, -24),
        to_sfixed(1.5258789061315762e-05, 7, -24),
        to_sfixed(7.62939453110197e-06, 7, -24),
        to_sfixed(3.814697265606496e-06, 7, -24),
        to_sfixed(1.907348632810187e-06, 7, -24),
        to_sfixed(9.536743164059608e-07, 7, -24),
        to_sfixed(4.7683715820308884e-07, 7, -24),
        to_sfixed(2.3841857910155797e-07, 7, -24),
        to_sfixed(1.1920928955078068e-07, 7, -24),
        to_sfixed(5.960464477539055e-08, 7, -24),
        to_sfixed(2.9802322387695303e-08, 7, -24),
        to_sfixed(1.4901161193847655e-08, 7, -24),
        to_sfixed(7.450580596923828e-09, 7, -24),
        to_sfixed(3.725290298461914e-09, 7, -24),
        to_sfixed(1.862645149230957e-09, 7, -24),
        to_sfixed(9.313225746154785e-10, 7, -24),
        to_sfixed(4.656612873077393e-10, 7, -24)
    );

    CONSTANT C_TANGENT_K32_CORR_TABLE_SFIXED: t_tan_ceoffs_sfixed(0 to 31) := (
        to_sfixed(0.4769353398736855, 7, -24),
        to_sfixed(0.4636476090008061, 7, -24),
        to_sfixed(0.24497866312686414, 7, -24),
        to_sfixed(0.12435499454676144, 7, -24),
        to_sfixed(0.06241880999595735, 7, -24),
        to_sfixed(0.031239833430268277, 7, -24),
        to_sfixed(0.015623728620476831, 7, -24),
        to_sfixed(0.007812341060101111, 7, -24),
        to_sfixed(0.0039062301319669718, 7, -24),
        to_sfixed(0.0019531225164788188, 7, -24),
        to_sfixed(0.0009765621895593195, 7, -24),
        to_sfixed(0.0004882812111948983, 7, -24),
        to_sfixed(0.00024414062014936177, 7, -24),
        to_sfixed(0.00012207031189367021, 7, -24),
        to_sfixed(6.103515617420877e-05, 7, -24),
        to_sfixed(3.0517578115526096e-05, 7, -24),
        to_sfixed(1.5258789061315762e-05, 7, -24),
        to_sfixed(7.62939453110197e-06, 7, -24),
        to_sfixed(3.814697265606496e-06, 7, -24),
        to_sfixed(1.907348632810187e-06, 7, -24),
        to_sfixed(9.536743164059608e-07, 7, -24),
        to_sfixed(4.7683715820308884e-07, 7, -24),
        to_sfixed(2.3841857910155797e-07, 7, -24),
        to_sfixed(1.1920928955078068e-07, 7, -24),
        to_sfixed(5.960464477539055e-08, 7, -24),
        to_sfixed(2.9802322387695303e-08, 7, -24),
        to_sfixed(1.4901161193847655e-08, 7, -24),
        to_sfixed(7.450580596923828e-09, 7, -24),
        to_sfixed(3.725290298461914e-09, 7, -24),
        to_sfixed(1.862645149230957e-09, 7, -24),
        to_sfixed(9.313225746154785e-10, 7, -24),
        to_sfixed(4.656612873077393e-10, 7, -24)
    );

END PACKAGE cordic_pkg;
