--==========================================================================================
-- This VVC was generated with Bitvis VVC Generator
--==========================================================================================


context vvc_context is
  library bitvis_vip_apb;
  use bitvis_vip_apb.vvc_methods_pkg.all;
  use bitvis_vip_apb.td_vvc_framework_common_methods_pkg.all;
  use bitvis_vip_apb.apb_bfm_pkg.t_apb_if;
  use bitvis_vip_apb.apb_bfm_pkg.t_apb_bfm_config;
  use bitvis_vip_apb.apb_bfm_pkg.C_APB_BFM_CONFIG_DEFAULT;
end context;
